module LCD_Display(iCLK_50MHZ, iRST_N, hex1, hex0, 
    LCD_RS,LCD_E,LCD_RW,DATA_BUS,botao, led0, led1, led2, led3,botao0,botao1,botao2, chave4);
input iCLK_50MHZ, iRST_N;
input [3:0] hex1, hex0;
output LCD_RS, LCD_E, LCD_RW;
inout [7:0] DATA_BUS;
input botao;
output led0,led1, led2, led3;
input botao0,botao1,botao2;
input [0:3]chave4;//Escolher produto

parameter
HOLD = 4'h0,
FUNC_SET = 4'h1,
DISPLAY_ON = 4'h2,
MODE_SET = 4'h3,
Print_String = 4'h4,
LINE2 = 4'h5,
RETURN_HOME = 4'h6,
DROP_LCD_E = 4'h7,
RESET1 = 4'h8,
RESET2 = 4'h9,
RESET3 = 4'ha,
DISPLAY_OFF = 4'hb,
DISPLAY_CLEAR = 4'hc;

reg [3:0] state, next_command;
// Enter new ASCII hex data above for LCD Display
reg [7:0] DATA_BUS_VALUE;
wire [7:0] Next_Char;
reg [19:0] CLK_COUNT_400HZ;
reg [4:0] CHAR_COUNT;
reg CLK_400HZ, LCD_RW_INT, LCD_E, LCD_RS;

// BIDIRECTIONAL TRI STATE LCD DATA BUS
assign DATA_BUS = (LCD_RW_INT? 8'bZZZZZZZZ: DATA_BUS_VALUE);

Maquina u1(
.index(CHAR_COUNT),
.out(Next_Char),
.hex1(hex1),
.hex0(hex0),
.botao(botao),
.led0(led0),
.led1(led1),
.led2(led2),
.led3(led3),
.clock(iCLK_50MHZ),
.botao0(botao0),
.botao1(botao1),
.botao2(botao2),
.chave4(chave4)
);

assign LCD_RW = LCD_RW_INT;

always @(posedge iCLK_50MHZ or negedge iRST_N)
    if (!iRST_N)
    begin
       CLK_COUNT_400HZ <= 20'h00000;
       CLK_400HZ <= 1'b0;
    end
    else if (CLK_COUNT_400HZ < 20'h0F424)
    begin
       CLK_COUNT_400HZ <= CLK_COUNT_400HZ + 1'b1;
    end
    else
    begin
      CLK_COUNT_400HZ <= 20'h00000;
      CLK_400HZ <= ~CLK_400HZ;
    end
// State Machine to send commands and data to LCD DISPLAY

always @(posedge CLK_400HZ or negedge iRST_N)
    if (!iRST_N)
    begin
     state <= RESET1;
    end
    else
    case (state)
    RESET1:            
// Set Function to 8-bit transfer and 2 line display with 5x8 Font size
// see Hitachi HD44780 family data sheet for LCD command and timing details
    begin
      LCD_E <= 1'b1;
      LCD_RS <= 1'b0;
      LCD_RW_INT <= 1'b0;
      DATA_BUS_VALUE <= 8'h38;
      state <= DROP_LCD_E;
      next_command <= RESET2;
      CHAR_COUNT <= 5'b00000;
    end
    RESET2:
    begin
      LCD_E <= 1'b1;
      LCD_RS <= 1'b0;
      LCD_RW_INT <= 1'b0;
      DATA_BUS_VALUE <= 8'h38;
      state <= DROP_LCD_E;
      next_command <= RESET3;
    end
    RESET3:
    begin
      LCD_E <= 1'b1;
      LCD_RS <= 1'b0;
      LCD_RW_INT <= 1'b0;
      DATA_BUS_VALUE <= 8'h38;
      state <= DROP_LCD_E;
      next_command <= FUNC_SET;
    end
// EXTRA STATES ABOVE ARE NEEDED FOR RELIABLE PUSHBUTTON RESET OF LCD

    FUNC_SET:
    begin
      LCD_E <= 1'b1;
      LCD_RS <= 1'b0;
      LCD_RW_INT <= 1'b0;
      DATA_BUS_VALUE <= 8'h38;
      state <= DROP_LCD_E;
      next_command <= DISPLAY_OFF;
    end

// Turn off Display and Turn off cursor
    DISPLAY_OFF:
    begin
      LCD_E <= 1'b1;
      LCD_RS <= 1'b0;
      LCD_RW_INT <= 1'b0;
      DATA_BUS_VALUE <= 8'h08;
      state <= DROP_LCD_E;
      next_command <= DISPLAY_CLEAR;
    end

// Clear Display and Turn off cursor
    DISPLAY_CLEAR:
    begin
      LCD_E <= 1'b1;
      LCD_RS <= 1'b0;
      LCD_RW_INT <= 1'b0;
      DATA_BUS_VALUE <= 8'h01;
      state <= DROP_LCD_E;
      next_command <= DISPLAY_ON;
    end

// Turn on Display and Turn off cursor
    DISPLAY_ON:
    begin
      LCD_E <= 1'b1;
      LCD_RS <= 1'b0;
      LCD_RW_INT <= 1'b0;
      DATA_BUS_VALUE <= 8'h0C;
      state <= DROP_LCD_E;
      next_command <= MODE_SET;
    end

// Set write mode to auto increment address and move cursor to the right
    MODE_SET:
    begin
      LCD_E <= 1'b1;
      LCD_RS <= 1'b0;
      LCD_RW_INT <= 1'b0;
      DATA_BUS_VALUE <= 8'h06;
      state <= DROP_LCD_E;
      next_command <= Print_String;
    end

// Write ASCII hex character in first LCD character location
    Print_String:
    begin
      state <= DROP_LCD_E;
      LCD_E <= 1'b1;
      LCD_RS <= 1'b1;
      LCD_RW_INT <= 1'b0;
    // ASCII character to output
      if (Next_Char[7:4] != 4'h0)
        DATA_BUS_VALUE <= Next_Char;
        // Convert 4-bit value to an ASCII hex digit
      else if (Next_Char[3:0] >9)
        // ASCII A...F
         DATA_BUS_VALUE <= {4'h4,Next_Char[3:0]-4'h9};
      else
        // ASCII 0...9
         DATA_BUS_VALUE <= {4'h3,Next_Char[3:0]};
    // Loop to send out 32 characters to LCD Display  (16 by 2 lines)
      if ((CHAR_COUNT < 31) && (Next_Char != 8'hFE))
         CHAR_COUNT <= CHAR_COUNT + 1'b1;
      else
         CHAR_COUNT <= 5'b00000; 
    // Jump to second line?
      if (CHAR_COUNT == 15)
        next_command <= LINE2;
    // Return to first line?
      else if ((CHAR_COUNT == 31) || (Next_Char == 8'hFE))
        next_command <= RETURN_HOME;
      else
        next_command <= Print_String;
    end

// Set write address to line 2 character 1
    LINE2:
    begin
      LCD_E <= 1'b1;
      LCD_RS <= 1'b0;
      LCD_RW_INT <= 1'b0;
      DATA_BUS_VALUE <= 8'hC0;
      state <= DROP_LCD_E;
      next_command <= Print_String;
    end

// Return write address to first character postion on line 1
    RETURN_HOME:
    begin
      LCD_E <= 1'b1;
      LCD_RS <= 1'b0;
      LCD_RW_INT <= 1'b0;
      DATA_BUS_VALUE <= 8'h80;
      state <= DROP_LCD_E;
      next_command <= Print_String;
    end

// The next three states occur at the end of each command or data transfer to the LCD
// Drop LCD E line - falling edge loads inst/data to LCD controller
    DROP_LCD_E:
    begin
      LCD_E <= 1'b0;
      state <= HOLD;
    end
// Hold LCD inst/data valid after falling edge of E line                
    HOLD:
    begin
      state <= next_command;
    end
    endcase
endmodule

module Maquina(index,out,hex0,hex1,clock, botao0,botao1,botao2,chave4, led0, led1, led2, led3,botao);
input [4:0] index;
input [3:0] hex0,hex1;
output [7:0] out;
reg [7:0] out;
input clock, botao;
input botao0,botao1,botao2; //Receber o dinheiro
input [0:3]chave4;//Escolher produto
output led0, led1, led2, led3;
reg [3:0] soma, totalAPagar,troco;
reg estadoLed0, estadoLed1, estadoLed2, estadoLed3;
reg [1:0] estado;
reg[31:0] contador, contador1; // REGISTRA 32 DIGITOS
wire chave0,chave1,chave2,chave3;

initial begin
contador <= 32'b0;// ZERA O CONTADOR
contador1 <= 32'b0;// ZERA O CONTADOR
soma <= 0;// ZERA O CONTADOR
totalAPagar <= 0;// ZERA O CONTADOR
troco <= 0;
end

parameter zero=0, um=1, dois=2, tres=3;

always @(posedge clock) 
begin
	case (estado)
		zero:
			begin
			estadoLed0 <= 1'b1;
			estadoLed1 <= 1'b0;
			estadoLed2 <= 1'b0;
			estadoLed3 <= 1'b0;
			
			case (index)
								5'h00: out <= 8'h53; //s
								5'h01: out <= 8'h65; //e
								5'h02: out <= 8'h6C; //l
								5'h03: out <= 8'h65; //e
								5'h04: out <= 8'h63; //c
								5'h05: out <= 8'h69; //i
								5'h06: out <= 8'h6F; //o
								5'h07: out <= 8'h6E; //n
								5'h08: out <= 8'h65; //e
								5'h09: out <= 8'h20; //espaco
								5'h0A: out <= 8'h56; //v
								5'h0B: out <= 8'h61; //a
								5'h0C: out <= 8'h6C; //l
								5'h0D: out <= 8'h6F; //o
								5'h0E: out <= 8'h72; //r
								
								// Line 2
								5'h10: out <= 8'h56; //v
								5'h11: out <= 8'h61; //a
								5'h12: out <= 8'h6C; //l
								5'h13: out <= 8'h6F; //o
								5'h14: out <= 8'h72; //r
								default: out <= 8'h20;
			endcase
			if(~botao0 || ~botao1 || ~botao2)
			begin
			contador1 <= contador1 + 1'b1; // SOMA UM AO CONTADOR
			end
			
			if(contador1 > 15000000) // SE O CONTADOR = MÁXIMO
			begin
				if(~botao0)
				begin
				soma <= soma + 4'b0001; // SOMA UM 
				end
				if(~botao1)
				begin
				soma <= soma + 4'b0010; // SOMA UM 
				end
				if(~botao2)
				begin
				soma <= soma + 4'b0101;
				end
				contador1 <= 0; // ZERA CONTADOR
			end
			
			case (soma)
			4'b0000:
			begin
			case (index)
				5'h15: out <= 8'h20; //espaco
				5'h16: out <= 8'h30;
			endcase
			end //espaco
			4'b0001:
			begin
			case (index)
				5'h15: out <= 8'h20; //espaco
				5'h16: out <= 8'h31;
			endcase
			end //espaco
			4'b0010:
			begin
			case (index)
				5'h15: out <= 8'h20; //espaco
				5'h16: out <= 8'h32; //espaco
			endcase
			end
			4'b0011:
			begin
			case (index)
				5'h15: out <= 8'h20; //espaco
				5'h16: out <= 8'h33; //espaco
			endcase
			end
			4'b0100:
			begin
			case (index)
				5'h15: out <= 8'h20; //espaco
				5'h16: out <= 8'h34; //espaco
			endcase
			end
			4'b0101:
			begin
			case (index)
				5'h15: out <= 8'h20;//espaco
				5'h16: out <= 8'h35; //espac
			endcase
			end
			4'b0110:
			begin
			case (index)
				5'h15: out <= 8'h20; //espaco
				5'h16: out <= 8'h36; //espaco
			endcase
			end
			4'b0111:
			begin
			case (index)
				5'h15: out <= 8'h20; //espaco
				5'h16: out <= 8'h37; //espaco
			endcase
			end
			4'b1000:
			begin
			case (index)
				5'h15: out <= 8'h20; //espaco
				5'h16: out <= 8'h38; //espaco
			endcase
			end
			endcase
			
			
	end
		um:
			begin
			estadoLed0 <= 1'b0;
			estadoLed1 <= 1'b1;
			estadoLed2 <= 1'b0;
			estadoLed3 <= 1'b0; 
			
			case (index)
							5'h00: out <= 8'h53; //s
							5'h01: out <= 8'h65; //e
							5'h02: out <= 8'h6C; //l
							5'h03: out <= 8'h65; //e
							5'h04: out <= 8'h63; //c
							5'h05: out <= 8'h69; //i
							5'h06: out <= 8'h6F; //o
							5'h07: out <= 8'h6E; //n
							5'h08: out <= 8'h65; //e
							// Line 2
							5'h10: out <= 8'h6F; //o
							5'h11: out <= 8'h20; //espaco
							5'h12: out <= 8'h70; //p
							5'h13: out <= 8'h72; //r
							5'h14: out <= 8'h6F; //o
							5'h15: out <= 8'h64; //d
							5'h16: out <= 8'h75; //u
							5'h17: out <= 8'h74; //t
							5'h18: out <= 8'h6F; //o
							5'h19: out <= 8'h3A; //:
							default: out <= 8'h20;
			endcase
			case(chave4)
					4'b0000:
						totalAPagar = 4'b0000;
					4'b0001:
						totalAPagar = 4'b0010;
					4'b0010:
						totalAPagar = 4'b0010;
					4'b0011:
						totalAPagar = 4'b0100;
					4'b0100:
						totalAPagar = 4'b0010;
					4'b0101:
						totalAPagar = 4'b0100;
					4'b0110:
						totalAPagar = 4'b0100;
					4'b0111:
						totalAPagar = 4'b0110;
					4'b1000:
						totalAPagar = 4'b0010;
					4'b1001:
						totalAPagar = 4'b0100;
					4'b1010:
						totalAPagar = 4'b0100;
					4'b1011:
						totalAPagar = 4'b0110;
					4'b1100:
						totalAPagar = 4'b0100;
					4'b1101:
						totalAPagar = 4'b0110;
					4'b1110:
						totalAPagar = 4'b0110;
					4'b1111:
						totalAPagar = 4'b1000;
				endcase
			end
		dois:
			begin
			estadoLed0 <= 1'b0;
			estadoLed1 <= 1'b0;
			estadoLed2 <= 1'b1;
			estadoLed3 <= 1'b0;
			
			case (index)     		
								5'h00: out <= 8'h70; //p
								5'h01: out <= 8'h72; //r
								5'h02: out <= 8'h6F; //o
								5'h03: out <= 8'h64; //d
								5'h04: out <= 8'h75; //u
								5'h05: out <= 8'h74; //t
								5'h06: out <= 8'h6F; //o
								5'h07: out <= 8'h20; //espaco
								5'h08: out <= 8'h73; //s
								5'h09: out <= 8'h61; //a
								5'h0a: out <= 8'h69;//i
								5'h0b: out <= 8'h6E;//n
								5'h0c: out <= 8'h64;//d
								5'h0d: out <= 8'h6F;//o
								// Line 2
								5'h10: out <= 8'h74; //t
								5'h11: out <= 8'h72; //r
								5'h12: out <= 8'h6F; //o
								5'h13: out <= 8'h63; //c
								5'h14: out <= 8'h6F; //o
								5'h15: out <= 8'h20; //espaco
								5'h16: out <= 8'h3D; //=
								5'h17: out <= 8'h20; //espaco
								default: out <= 8'h20;
								
								
			endcase
			troco = totalAPagar - soma;
			case (troco)
				4'b0000:
				begin
				case (index)
					5'h18: out <= 8'h30;
				endcase
				end //espaco
				4'b0001:
				begin
				case (index)
					5'h18: out <= 8'h31;
				endcase
				end //espaco
				4'b0010:
				begin
				case (index)
					5'h18: out <= 8'h32; //espaco
				endcase
				end
				4'b0011:
				begin
				case (index)
					5'h18: out <= 8'h33; //espaco
				endcase
				end
				4'b0100:
				begin
				case (index)
					5'h18: out <= 8'h34; //espaco
				endcase
				end
				4'b0101:
				begin
				case (index)
					5'h18: out <= 8'h35; //espac
				endcase
				end
				4'b0110:
				begin
				case (index)
					5'h18: out <= 8'h36; //espaco
				endcase
				end
				4'b0111:
				begin
				case (index)
					5'h18: out <= 8'h37; //espaco
				endcase
				end
				4'b1000:
				begin
				case (index)
					5'h18: out <= 8'h38; //espaco
				endcase
				end
			endcase

			end
		tres:
			begin
			estadoLed0 <= 1'b0;
			estadoLed1 <= 1'b0;
			estadoLed2 <= 1'b0;
			estadoLed3 <= 1'b1;
			
			case (index)
								5'h00: out <= 8'h74; //t
								5'h01: out <= 8'h65; //e
								5'h02: out <= 8'h6E; //n
								5'h03: out <= 8'h74; //t
								5'h04: out <= 8'h61; //a
								5'h05: out <= 8'h72; //r
								5'h06: out <= 8'h20; //espaco
								// Line 2
								5'h10: out <= 8'h6E; //n
								5'h11: out <= 8'h6F; //o
								5'h12: out <= 8'h76; //v
								5'h13: out <= 8'h61; //a
								5'h14: out <= 8'h6D; //m
								5'h15: out <= 8'h65; //e
								5'h16: out <= 8'h6E; //n
								5'h17: out <= 8'h74; //t
								5'h18: out <= 8'h65; //e
								default: out <= 8'h20;
			endcase
			end
		default:
			begin
			estadoLed0 <= 1'b0;
			estadoLed1 <= 1'b0;
			estadoLed2 <= 1'b0;
			estadoLed3 <= 1'b0;
			end
	endcase
end

always @(posedge clock) // SEMPRE NO PULSO DO CLOCK
begin
	if(~botao)
	begin
	contador <= contador + 1'b1; // SOMA UM AO CONTADOR
	end
	
	if(contador > 15000000) // SE O CONTADOR = M�XIMO
	begin
		case (estado)
			zero:
				 estado = um;
			um:
				 if(soma >= totalAPagar && totalAPagar>0)
					estado = dois;
				 else
					estado = tres;
			dois:
				estado = zero;
			tres:
				estado = zero;
        endcase
		contador <= 0; // ZERA CONTADOR
	end
end

assign led0 = estadoLed0; // LED � ASSOCIADO AO ESTADO
assign led1 = estadoLed1; // LED � ASSOCIADO AO ESTADO
assign led2 = estadoLed2; // LED � ASSOCIADO AO ESTADO
assign led3 = estadoLed3; // LED � ASSOCIADO AO ESTADO

endmodule


